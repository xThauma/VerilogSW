module PS2_ZAD9(
	output [6:0] HEX0, HEX1, HEX2, HEX3);

		assign HEX0=7'b0100011;		//	o
		assign HEX1=7'b0000111;		// t
		assign HEX2=7'b1100011;		// u
		assign HEX3=7'b0100000;		// a

endmodule
