module PS2_ZAD10(
	output [6:0] HEX0, HEX1, HEX2, HEX3, HEX4, HEX5);
		assign HEX0=7'b0100011;		//	o
		assign HEX1=7'b0000111;		// t
		assign HEX2=7'b1111111; 	//spacja
		assign HEX3=7'b1111111; 	//spacja
		assign HEX4=7'b1100011;		// u
		assign HEX5=7'b0100000;		// a
		
endmodule
